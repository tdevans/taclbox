library ieee;
use ieee.std_logic_1164.all;

package types is
	type t_slv_array is array (natural range <>) of std_logic_vector;
end package types;